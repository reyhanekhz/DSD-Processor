module control_unit (
    input clk, reset, start,
    output reg ready,
    output reg [9:0] mem_address,
    output reg mem_write_enable, mem_read_enable,
    output reg signed [15:0] mem_data_in,
    input signed [15:0] mem_data_out,
    output reg reg_write_enable,
    output reg [1:0] reg_read_addr1, reg_read_addr2, reg_write_addr,
    output reg signed [15:0] reg_write_data,
    input signed [15:0] reg_read_data1, reg_read_data2,
    output reg alu_start,
    output reg [2:0] alu_opcode,
    output reg signed [15:0] alu_a, alu_b,
    input signed [15:0] alu_result_low, alu_result_high,
    input alu_done
);

    // States
    parameter IDLE          = 4'd0;
    parameter FETCH         = 4'd1;
    parameter ACCESS_MEMORY = 4'd2;
    parameter DECODE        = 4'd3;
    parameter EXECUTE       = 4'd4;
    parameter RF_ACCESS     = 4'd5;
    parameter ALU_WAIT      = 4'd6;
    parameter MEMORY        = 4'd7;
    parameter WRITEBACK     = 4'd8;
    parameter COMPLETE      = 4'd9;
    reg [3:0] state, previous_state;



    // PC register
    reg [9:0] PC;

    reg [15:0] instr;
    reg [2:0] opcode;
    reg [1:0] rd, rs1, rs2, base;
    reg [8:0] address_imm;       

    reg [9:0] effective_addr; // Address for load/store




    always @(posedge clk or posedge reset) begin
        // Reset everything and set state as IDLE in the beginning
        if (reset) begin
            PC <= 10'b0;
            state <= IDLE;
            ready <= 1'b0;
            mem_read_enable <= 1'b0;
            mem_write_enable <= 1'b0;
            reg_write_enable <= 1'b0;
            alu_start <= 1'b0;
        end 
        
        else begin
            case (state)
                IDLE: begin
                    ready <= 0;
                    if (start) begin
                        state <= FETCH;
                        previous_state <= IDLE;
                    end
                end

                FETCH: begin // read instruction from memory 
                    mem_address <= PC;
                    mem_read_enable <= 1'b1;
                    ready <= 1'b0;
                    state <= ACCESS_MEMORY;
                    previous_state <= FETCH;
                end

                ACCESS_MEMORY: begin // One cycle to read form memory
                    mem_read_enable <= 1'b0;

                    // Writeback to register file when LOAD
                    if (previous_state == MEMORY) begin
                        state <= WRITEBACK;
                        previous_state <= ACCESS_MEMORY;
                    end

                    else begin
                        state <= DECODE;
                        previous_state <= ACCESS_MEMORY;
                    end
                end

                DECODE: begin
                    instr <= mem_data_out;

                    opcode <= mem_data_out[15:13];

                    // M-type format
                    if (mem_data_out[15:13] == 3'b100 || mem_data_out[15:13] == 3'b101) begin
                        rd <= mem_data_out[12:11];
                        base <= mem_data_out[10:9];
                        address_imm <= mem_data_out[8:0];
                        state <= EXECUTE;
                        previous_state <= DECODE;
                    end 
                    
                    // R-type format
                    else begin
                        rd <= mem_data_out[12:11];
                        rs1 <= mem_data_out[10:9];
                        rs2 <= mem_data_out[8:7];
                        state <= EXECUTE;
                        previous_state <= DECODE;
                    end
                end

                EXECUTE: begin
                    if (opcode == 3'b100 || opcode == 3'b101) begin
                        reg_read_addr1 <= base;
                        // Read rd to store in memory
                        if (opcode == 3'b101) begin
                            reg_read_addr2 <= rd;
                        end
                        state <= RF_ACCESS;
                        previous_state <= EXECUTE;
                    end 
                    
                    else begin
                        reg_read_addr1 <= rs1;
                        reg_read_addr2 <= rs2;
                        state <= RF_ACCESS;
                        previous_state <= EXECUTE;
                    end
                end

                RF_ACCESS: begin // One half-cycle to access register file
                    if (opcode == 3'b100 || opcode == 3'b101) begin
                        effective_addr <= reg_read_data1[9:0] + {address_imm[8], address_imm};
                        state <= MEMORY;
                        previous_state <= RF_ACCESS;
                    end

                    else begin
                        alu_a <= reg_read_data1;
                        alu_b <= reg_read_data2;
                        alu_opcode <= opcode;
                        alu_start <= 1'b1;

                        state <= ALU_WAIT;
                        previous_state <= RF_ACCESS;
                    end
                end

                ALU_WAIT: begin
                    // Wait till ALU is done
                    if (alu_done) begin
                        alu_start <= 1'b0;
                        reg_write_addr <= rd;
                        reg_write_data <= alu_result_low[15:0];
                        reg_write_enable <= 1'b1;
                        state <= WRITEBACK;
                        previous_state <= ALU_WAIT;
                    end
                end

                MEMORY: begin
                    // Load
                    if (opcode == 3'b100) begin
                        mem_address <= effective_addr;
                        mem_read_enable <= 1'b1;
                        state <= ACCESS_MEMORY;
                        previous_state <= MEMORY;
                    end 
                    
                    // Store
                    else begin
                        mem_address <= effective_addr;
                        mem_write_enable <= 1'b1;
                        mem_data_in <= reg_read_data2;
                        state <= COMPLETE;
                        previous_state <= MEMORY;
                    end
                end
 
                WRITEBACK: begin
                    mem_read_enable <= 1'b0;
                    if (opcode == 3'b100) begin
                        reg_write_enable <= 1'b1;
                        reg_write_addr <= rd;
                        reg_write_data <= mem_data_out;
                    end
                    state <= COMPLETE;
                    previous_state <= WRITEBACK;
                end

                COMPLETE: begin
                    reg_write_enable <= 1'b0;
                    mem_write_enable <= 1'b0;
                    alu_start <= 1'b0;
                    PC <= PC + 1;
                    ready <= 1'b1;
                    state <= FETCH;
                    previous_state <= COMPLETE;
                end

            endcase
        end
    end
endmodule
